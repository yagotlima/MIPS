LIBRARY	ieee;
USE		ieee.std_logic_1164.all;

entity MIPS is
	port(
		CLK, RESET	: in  STD_LOGIC;
	);
end MIPS;

architecture mips_arch of MIPS is
begin
	-- TODO --
end;
